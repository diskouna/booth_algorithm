package utils is 
    function clog2(number : positive) return positive;
end package;

package body utils is
    function clog2(number : positive) return positive is
        variable numbers_bits : positive := 8;
    begin 
        --TODO       
        return numbers_bits;
    end function;
end package body;
